program testcase();
 //import uvm_pkg::*;

 //`include "../../testbench/verilog_new/uvm_test_top.sv"

  initial begin
    run_test("uvm_test_top");
  end	
endprogram  


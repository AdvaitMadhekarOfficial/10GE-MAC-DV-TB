interface reset_if(input wb_clk_i, input clk_156m25);
  logic wb_rst_i;
  logic reset_156m25_n;
endinterface
